library ieee;
use ieee.std_logic_1164.all;

entity Test_RegistroUniversal is
end  Test_RegistroUniversal;
